module adder(a, b, out);
input [63:0] a, b;
output [63:0] out;
assign out = a + b;
endmodule;1
