module program_counter(in,out);
input [63:0] in;
output reg [63:0] out;

always
begin
out=in;
end
endmodule;1
